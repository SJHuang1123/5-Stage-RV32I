module imem_1024x32(
  input  [9:0]  R0_addr,
  input         R0_en,
                R0_clk,
  output [31:0] R0_data
);

  reg [31:0] Memory[0:1023];
  assign R0_data = R0_en ? Memory[R0_addr] : 32'bx;
endmodule

module InstMem(
  input         clock,
                reset,
  input  [31:0] io_addr,
  output [31:0] io_data
);

  wire [31:0] _io_data_T = io_addr / 32'h4;
  imem_1024x32 imem_ext (
    .R0_addr (_io_data_T[9:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R0_data (io_data)
  );
endmodule
// ----- 8< ----- FILE "imem_1024x32_init.sv" ----- 8< -----

// Generated by CIRCT firtool-1.62.1
module imem_1024x32_init();
  initial
    $readmemh("test.txt", imem_1024x32.Memory);
endmodule

bind imem_1024x32 imem_1024x32_init imem_1024x32_init ();
